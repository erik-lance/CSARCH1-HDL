//Test bench
`include "tioe1.v"

module tioe1_tb;


endmodule