//test
module tioe1(A, B, C, D);



endmodule